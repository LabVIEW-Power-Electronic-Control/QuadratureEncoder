-- � 2012 National Instruments Corporation.
encrypted

�U��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D���[�
d�U���u�0�0�4�2�}�ψ�����g+�"��Xʝ�2�x�0�0�w�$�����ƪ�\��N��^ʴ�1��&�0��p�W���
����T��@�X���:�,�<�=�w��W��MӾ��Z��~ ��U���u�<�=�&�%�.����W���9K�
S��H��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D����Z��E��0���_�&�u���.��������P��V�����u���;�:�/����݇��l��Y��ʸ�f�����}������F�V�����u������4�ԜY�ƭ�l��T��;ʆ�����]�}�W���
����\��yN��1�����_�u�w�-����Y�ƃ�gF��s1��2���_�u�u�%�>�1�W���,�Ɵ�w9��p'�����u�%�'�4�.�g�8���*����|!��d��Uʥ�e��1�0��>�Mϑ�-ӵ��l*��~-��0����}�d�1� �)�W���s���C9��e�����6�4�
�9�w�}�"���-����t/��=N��U���
�=�!�u�w��W���&����p9��t:��U��u�:�;�:�g�f�W���	�ד�[��h�����o������0���s���C9��e�����6�o�����;���:����g)��]����!�u�|�_�w�}�(݁�����`��V�����u� �u����>��Y����lU��R�� ���;�u�u� �w�	�(���0����p2��F�U���;�:�e�n�w�}����+����F��Y�����1�o�����;���:���F��1��%���0�u�u����;���:����g)��]����!�u�|�_�w�}����Y�ƅ�5��h"��<��u�u�%�c�3�����&����_�'��&������_�w�}�(ׁ�����c��RN�<����
�����#���Q����\��XN�N���u�%�m��!�8�'�������E
��N��U���
���n�w�}���&����\��^��Oʜ�u��
����2���+������Y��E��u�u�%�d��8�'�������R��[
��U��������W�W���&�ד�Q��D�����u������4���:����U��S�����|�_�u�u��l�6�������\��G1�����u��
���W������9l��T�����'�u�0�4�w�;���;����U9��^��U���4�!�<� �2��%���<����g/��h'��:�����n�w�}��������%��r1��;�����
���2�W�������R��^�����u�&�u�u�u�m�E���=������h��G��
�y�����#���)�ۯ�KJ��d1��%������d���>���-����v"�&��*��� �
���/�j�G�������W��{=��;���
���h�b�m�G��U����z(��c1��6���!�0�&����9���6���H��^�Y���
��
��j�m�?���*����c2��X ��=�������g��$���7����^��{=��,����d�m�y���.���,����R��d��Uʶ�;�!�;�u�'�>��������lW�=��*����u�h�r�p�W�W�������]��G1�����9�2�6�e�m��3���>���F�UךU���:�&�4�!�6��#���H����lV�=��*����
����u�GϺ�����O�
N��E��e�e�e�w�]�}�W���
������d:��؊�&�
�u�u���8���&����|4�^�����:�e�u�h�u�m�G��I����l�N�����;�u�%���)�(���&����`2��{!��6�����u�d�w�2����I����D��^�E��e�n�u�u�4�3����Y����g9��1����o������!���6���F��@ ��U���o�u�e�e�g�m�G��B�����D��ʴ�
��&�`�1�0�C��*����|!��h8��!���}�e�1�"�#�}�^��Y����V��^�W�ߊu�u�:�&�6�)����-����l ��h[��U���
���
��	�%���Iӂ��]��G��H���e�e�d�e�g��}���Y����G����&���!�
�&�
�w�}�#���6����e#��x<��D���:�;�:�e�w�`�U��I����V��d��Uʶ�;�!�;�u�'��(���&����F��d:��9�������w�l�W������F��L�E��e�e�e�n�w�}��������R��c1��L���8�m�o����0���/����aF�N�����u�|�o�u�g�l�G��I���9F������!�4�
��$�l�(���&����`2��{!��6�����u�d�w�2����I����D��^�E��e�n�u�u�4�3����Y����g9��_�����e�o�����4���:����W��S�����|�o�u�d�g�m�G��I��ƹF��X �����4�
�:�&��+�E��Cӵ��l*��~-��0����}�d�1� �)�W���C���V��^�E��e�e�e�e�g�m�G��I���9F������!�4�
�:�$��ށ�Y�Ɵ�w9��p'��#����u�e�1� �)�W���C���]ǻN�����4�!�4�
�8�.�(���K���5��h"��<������}�f�9� ���Y���F�^�E��e�e�e�e�g�m�G��I����W�=N��U���&�4�!�4��2�����ԓ�\��c*��:���
�����l��������\�^�E��e�e�e�e�g�m�G��I����V��UךU���:�&�4�!�6�����&����lU�=��*����
����u�FϺ�����O�
N��E��e�e�e�e�g�m�G��I����V��_�����u�:�&�4�#�<�(���
���� T��T��!�����
����_������\F��T��W��e�e�e�e�g�m�G��I����V��_�W�ߊu�u�:�&�6�)��������_��hY��U���
���
��	�%���Hӂ��]��G��H���e�e�e�e�g�m�G��I����V��^�D���_�u�u�:�$�<�Ͽ�&����G9��\��U����
�����#���Q����\��XN�U��w�e�e�e�g�m�G��I����V��^�D��w�_�u�u�8�.��������]��[�*���u��
����2���+������Y��E���h�w�e�e�g�m�G��I����V��^�E��e�w�_�u�w�2����Ӈ��P	��C1��F؊�u�u��
���(���-��� W��X����u�h�w�e�g�m�G��I����V��^�E��d�d�w�_�w�}��������C9��Y����
�e�e�e�g�g�$���5����l0��c!��]��1�"�!�u�~�g�W��I����V��^�E��e�e�e�e�g�m�G��Y����\��V �����:�&�
�#�e�i�G��I����`2��{!��6�����u�f�w�2����I����D��^�E��e�e�e�e�g�m�G��I����D��N�����!�;�u�%�4�3����J����	F��s1��2������u�d�}�������	[�^�E��e�e�e�e�g�m�G��I����V��d��Uʶ�;�!�;�u�'�>��������V��(��U����
�����#���Q����\��XN�U��w�d�e�e�g�l�G��H����W��_�D��w�_�u�u�8�.��������]��[�*ٓ�e�e�e�o���;���:����g)��]����!�u�|�o�w�m�F��H����V��^�E��e�e�e�e�g�f�W�������R��V�����
�#�g��o�m�G���Y����)��t1��6���u�f�u�:�9�2�G���D����W��_�E��e�e�e�e�g�m�G��I����F�T�����u�%�6�;�#�1�D݁�N����g"��x)��*�����}�d�3�*����P���V��^�E��e�e�e�e�g�m�G��H����]ǻN�����4�!�4�
�8�.�(���K�׉�	F��s1��2������u�d�}�������	[�^�E��e�e�e�e�g�m�G��I����W��d��Uʶ�;�!�;�u�'�>�����ޓ�\��c*��:���
�����}�������	[�^�E��w�_�u�u�8�.��������]��[�*���u��
����2���+������Y��E���h�w�e�e�g�m�G��I����V��L�U���6�;�!�;�w�-��������9��^��U���
���
��	�%���Mӂ��]��G��H���e�e�e�e�g�m�G���s���P	��C��U���6�;�!�9�f��C��Cӵ��l*��~-��0����}�a�1� �)�W���C���V��^�E��e�w�_�u�w�2����Ӈ��P	��C1��M���u�u��
���(���-���F��@ ��U���o�u�d�d�f�l�U�ԜY�Ư�]��Y�����;�!�9�d��m�W���-����t/��a+��:���d�u�:�;�8�m�W��[����V��^�E��n�u�u�6�9�)����	����@��A_��D��o������!���6���F��@ ��U���o�u�e�e�g�l�G��I���9F������!�4�
�:�$�����M���5��h"��<������}�c�9� ���Y���F�^�E��e�e�e�w�]�}�W���
������T�����d�
�u�u���8���&����|4�N�����u�|�o�u�g�m�G��I����F�T�����u�%�6�;�#�1�Fׁ�Y�Ɵ�w9��p'��#����u�d�u�8�3���Y���V��^�E��e�e�e�w�]�}�W���
������T�����d�
��o���;���:����g)��_����!�u�|�o�w�m�G��I����W��_�N���u�6�;�!�9�}��������ET��T��!�����
����_�������V�S��E���_�u�u�:�$�<�Ͽ�&����G9��1�Oʆ�������8���Iӂ��]��G��H���w�_�u�u�8�.��������]��[��D��������4���Y����\��XN�U��w�d�n�u�w�>�����ƭ�l��D�����`�o�����4���:����U��S�����|�o�u�e�g�m�G��I����V��^�E��e�d�d�n�w�}��������R��X ��*���
�u�u����>���<����N��S�����|�o�u�e�g�m�L���YӅ��@��CN��*���&�
�#�
�w�}�#���6����e#��x<��Aʱ�"�!�u�|�m�}�G��I��ƓF�D�����%��
�&�w�}�#���6����e#��x<��D���:�;�:�e�w�`�U��I����V��d��Uʴ�!�<� �0�1�0��������	F��E��N���u�4�!�<�"�8��������Z��X�����
�&�u�u�>�3�Ϸ�Yш��VD��N�����4�u�%�&�0�>����-����l ��h^��U���
���n�w�}�����ƭ�l��h��*��o�����W�W���������h
�����6�<�
�<�w�}�#���6����e#��x<��F���:�;�:�e�l�}�Wϭ�����C9��S:�����
�'�2�o���;���:����g)��]����!�u�|�o�w�m�G��I����V��^�E��e�e�e�e�g�f�W���
����_F��1��%���0�
�%�#�3�4�(���Y�Ɵ�w9��p'�����u�<�;�9�'�k��������R��[
�����o������M���I��ƹF��^	��ʥ�m��#�0��1����&����	F��s1��2������u�d�}�������9F������%�m��#�2�����	����	F��s1��2������u�d�}�������	[�^�E��e�e�e�e�g�m�G��I����V��d��Uʦ�2�4�u�
��8�'�������R��[
�����2�o�����4�ԜY�ƿ�T����*����'� �&��-����	����	F��s1��2���o�u�e�n�w�}�����Ƽ�V��R�����:�
�;�&�0�g�$���5����l0��c!��]��1�"�!�u�~�W�W���������1�����<�<�;�%�2�}�W���&����p9��t:��U��u�:�;�:�g�}�J���I����V��^�E��e�e�e�e�g�m�G���s���@��V��*����#�:�<�>�3��������l��T��!�����n�u�w�.����Y����l4��g�����
�%�#�1�'�8�W���-����t/��S��E��u�u�&�2�6�}�(���8����@��X �����2�o�����4���:����U��S�����|�_�u�u�>�3�Ϯ�H¹��@6��^�����0�u�u����>���<����N��
�����e�u�h�w�g�m�G��I����V��^�E��e�e�e�w�]�}�W�������lW��v�����<�;�4�
�;���������g"��x)��N���u�&�2�4�w��F���
����G��h�����%�0�u�u���8���Y���A��N�����4�u�����4�������W��T��!�����
����_������\F��T��W��e�e�e�e�g�m�G��I����V��^�W�ߊu�u�<�;�;�<�(���&����
S�,��9���n�u�u�&�0�<�W���&����U��N�&���������W��Y����G	�UךU���<�;�9�3��2��������9��P1�G��������4���Y����W	��C��\�ߊu�u�<�;�;�<�(���&����l5��D�����d�o�����4�ԜY�ƿ�T�������7�1�d�f�m��8���7���F��P ��U���
� �d�b�'�}�W���&����p9��t:��U��u�:�;�:�g�f�W���
����_F��h �����'�
�d�
�2��N���Y����)��t1��6���u�f�u�:�9�2�G��Y����Z��[N��*����g��!�e��(���J�ޓ� F��d:��9�������w�n�W������]ǻN�����9�3�
���o�8���Kʹ��A��^�Oʆ�������8���J�ƨ�D��^����u�<�;�9�0�-����L����\��c*��:���
�����l��������l�N�����u��-� �����&����V��N��1��������}�D�������V�=N��U���;�9�4�
�>�����*���� 9��Z1�Oʆ�����]�}�W�������C9��P1����b�o�����}���Y����R
��d1�� ����!�d�
�"�l�@���Y�Ɵ�w9��p'��#����u�f�u�8�3���B�����Y�������,� ��j����L���5��h"��<������}�f�9� ���Y����F�D�����:�9�-���)�D݁�����l��N��1��������}�GϺ�����O��N�����4�u�:�9�/�	�8���J����T9��N�&���������W������\F��d��Uʦ�2�4�u�%�$�:����&����GR��D��U����
���l�}�Wϭ�����R��^	�����f�u�u����L���Yӕ��]��V�����&�$��
�#�����Y�Ɵ�w9��p'�����u�<�;�9�6���������
F��u!��0���_�u�u�<�9�1����<����|��[��*���a�c�%�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����ƪ�l5��r-�� ���`�g�'�2�b�o�Mύ�=����z%��r-��'���d�1�"�!�w�t�}���Y����R
��X������!�f�
�"�i�@���Y�Ɵ�w9��p'��#����u�e�1� �)�W���s���@��V�����-���!�d�����M����`2��{!��6�����u�e�3�*����P���F��P ��U���&�2�6�0��	��������\��c*��:���n�u�u�&�0�<�W���
����W��_��U�����n�u�w�.����Y����U��Y��G��������4���Y����W	��C��\�ߊu�u�<�;�;�;�(���;����lT��E��@���o������!���6���F��@ ��U���_�u�u�<�9�1��������V��c1��L���8�m�o����0���s���@��V�����2�7�1�d�f�g�5���<����F�D������-� ���)�Eف�����F��d:��9�������w�n�W������]ǻN�����9�4�
�<��.����&����l ��hW��U���
���n�w�}�����ƭ�l��h��*��u�u����f�W���
����_F��h��*���$��
�!�f�;���Y�Ɵ�w9��p'�����u�<�;�9�6���������
F��u!��0���_�u�u�<�9�1��������9��T��!�����
����_������\F��d��Uʦ�2�4�u�'��(�F���	����`2��{!��6�����u�f�w�2����I��ƹF��^	��ʴ�
�<�
�&�&��(���&����F��d:��9����_�u�u�>�3�Ͽ�&����Q��^�Oʗ����_�w�}����Ӂ��l ��[�����u��
����2���+������Y��E��u�u�&�2�6�}��������l��N��1��������}�D�������V�=N��U���;�9�3�
������&�ѓ�F9�� 1��U����
�����#���Q����\��XN�N���u�&�2�4�w�����-����lW��Q��@݊�d�o�����4���:����U��S�����|�_�u�u�>�3�Ϲ�	����P��G^��U���
���
��	�%���Hӂ��]��G�U���&�2�4�u�%����N����	F��s1��2������u�d�}�������9F������2�%�3�
�`��G��*����|!��h8��!���}�d�1�"�#�}�^�ԜY�ƿ�T��	��*���d�d�%�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����Ƽ�e��h�� ��b�%�u�u���8���&����|4�_�����:�e�n�u�w�.����Y����e9��h_�*��o������!���6�����Y��E��u�u�&�2�6�}����&¹��lW��h�Oʆ�������8���K�ƨ�D��^����u�<�;�9�#�-�O�������V��G\��U���
���
��	�%���Y����G	�UךU���<�;�9�!�'�4����&����CT�=��*����
����u�W������]ǻN�����9�'�!�<�>�;�(��&���5��h"��<������}�c�9� ���Y����F�D�����8�
�
�
��(�E���	����`2��{!��6�����u�e�3�*����P���F��P ��U���
�8�d�3��n�(��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N�����%�
� �g�e�-�W���-����t/��a+��:���e�1�"�!�w�t�}���Y����R
��R��*���
�4�!�6�$����I����	F��s1��2������u�f�}�������9F������&�9�!�%�1��Eׁ�J����g"��x)��*�����}�a�3�*����P���F��P ��U���0� �!�&�1��Bف�J����g"��x)��*�����}�b�3�*����P���F��P ��U���-� ��;�"��N���&����e9��Q��Cފ�g�o�����4���:����W��S�����|�_�u�u�>�3�Ϫ�	�ӓ�F9��1��U����
�����#���Q�ƨ�D��^����u�<�;�9�#�-�A���&����CT�=��*����
����u�W������]ǻN�����9�!�%�3��e�(��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N�����3�
�l�
�d�g�$���5����l0��c!��]���:�;�:�e�l�}�Wϭ�����G��\�� ��a�%�u�u���8���&����|4� N�����u�|�_�u�w�4��������l ��^�����u��
����2���+����W	��C��\�ߊu�u�<�;�;�-�G��&¹��lT��h�Oʆ�������8���K�ƨ�D��^����u�<�;�9�#�-�F���&����CU�=��*����
����u�GϺ�����O��N�����4�u�
�0�"�)�C���&����CS�=��*����
����u�FϺ�����O��N�����4�u��-��	����&�ߓ�]9��c��*���g�m�%�u�w�	�(���0����p2��F�U���;�:�e�n�w�}�����ƿ�_9��GX�� ��e�%�u�u���8���&����|4�N�����u�|�_�u�w�4����
����^��Q��A܊�g�o�����4���:����V��X����n�u�u�&�0�<�W���&����l ��[�����u��
����2���+����W	��C��\�ߊu�u�<�;�;�;�(���5�Ԣ�F��1��*��
�d�o����0���/����aF�N�����u�|�_�u�w�4��������f*��x��D݊�:�<�!�3��k�(��Cӵ��l*��~-��0����}�d�1� �)�W���s���@��V�����
� �f�m�'�}�W���&����p9��t:��U��1�"�!�u�~�W�W���������h_�����b�
�d�o���;���:����g)��\����!�u�|�_�w�}����ӈ��A��Q��MҊ�g�o�����4���:����V��X����n�u�u�&�0�<�W�������F9��1��U����
�����#���Q�ƨ�D��^����u�<�;�9�#�-�C���&����CT�=��*����
����u�W������]ǻN�����9�2�%�3��j�(��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N��*����� �
�b�o��������lR��h�Oʆ�������8���J�ƨ�D��^����u�<�;�9�#�-�@���&����CR�=��*����
����u�W������]ǻN�����9�!�%�d��(�C���	����`2��{!��6�����u�g�w�2����I��ƹF��^	��ʻ�!�=�d�3��i�(��Cӵ��l*��~-��0����}�u�:�9�2�G��Y����Z��[N�����d�3�
�f��o�Mύ�=����z%��r-��'���u�:�;�:�g�f�W���
����_F��G1�*���a�d�%�u�w�	�(���0����p2��F����!�u�|�_�w�}����Ӂ��l ��Z�����1�u�u����>���<����N��S�����|�_�u�u�>�3�Ϲ�	����R��T��U���
���n�w�}�����ƭ�l��h�����
�!�
�&��}�W���&����p]ǻN�����9�4�
�<��9�(��Y�Ǝ�|*��yUךU���<�;�9�2�'�;�(��&���5��h"��<��u�u�&�2�6�}��������l��N��1�����_�u�w�4��������F9��1�����u�u��
���(���-���F��@ ��U���_�u�u�<�9�1����*����\��c*��:���
�����m��������l�N�����u�%�&�2�5�9�@���Y����v'��=N��U���;�9�4�
�>�����I����|)��v �U���&�2�4�u�'�.��������	F��x"��;�ߊu�u�<�;�;�<�(���&����T�,��9���n�_�u�u�8�-����Y����q'��v��*���1�&�7�f�9��E���J����U��h
��U���u�u�2�;�%�>�_���Y���/��N��!����_�u�u�w�}�"���-����	F��c+��'�ߊu�u�u�u�>�m� ���1����}2��r<�U���u�u�1�;���#���Y����t#��=N��U���u�:�!����Mϗ�-����O��N�����u�_�u�u�w�}����Y����g"��x)��N���u�u�u�'�$�)�Mϗ�Y����)��tUךU���u�u�<�e�m��W���&����p9��t:��U��u�:�;�:�g�f�W���Y����Z��N��U���
���
��	�%���Hӂ��]��G�U���u�u�:�6�3�}�W���*����|!��h8��!���}�u�:�;�8�m�L���Y�����N��U���
���n�w�}�W�������	F��cN��1��������}�D�������V�UךU���;�u�:�%�9�3�L�ԶY����\��Y��U��g���3�g�;����K������\��*���
�&�u��w�}�������9F�N��U���o�����W�W���Y�Ƃ�~9��v)��Oʜ����_�w�}�W����֓�z"��T��;����n�u�u�w�}����&����{F��~ ��2���_�u�u�u�w�2����=���/��r)��U��u�u�%�'�w�W�W���Y�ƨ�]V�'��&���������W��Y����G	�UךU���u�u�<�d�m��W���&����p9��t:��U��u�:�;�:�g�f�W���Y����\��N��!ʆ�������8���J�ƨ�D��^��\�ߊu�u�;�u�8�-����B��ƹF��X�����u�e�g���;�G������� T��h]��Gʜ�_�u�u�0�2�4�W�ԜY���F��T��;����n�u�u�w�}�9���*����\��y:��0��u�u�u�u�3�3�(���-����z(��p+�����u�u�u�:�#�
�3���Cӯ��v!��G�U���%�'�u�_�w�}�W�������z(��c*��:���n�u�u�u�w�/����Cӯ��`2��{!��6�ߊu�u�u�u�>�m�Mϗ�Y����)��t1��6���u�f�u�:�9�2�G��Y���F��RN�<����
���l�}�W���Yӂ��GF��x;��&���������W��Y����G	�N����u�;�u�:�'�3���s�����G�����e�g���1�m����&�Ԣ�lU��D1��Dʜ�_�u�u�0�2�4�W�ԜY���F��T��;����n�u�u�w�}�9���*����\��y:��0��u�u�u�u�3�3�(���-����z(��p+�����u�u�u�<�f�
�3���Cӯ��v!��d��U���u�1� �
��	�W���7����aF�=N��U���!�}�u�u�w�}����Y�ƅ�5��h"��<������}�f�9� ���Y����F�N�����u�u�����0���/����aF�N�����u�|�_�u�w�}�W������/��d:��9�������w�i��������l�N��Uʱ� �u�u� �w�	�(���0����p2��F����!�u�|�|�]�}�W���Y����\��CUװ��2�;�u�u�1�m�������� T��h]����
�
� �9�3�-�"���Y����\��CN��Fؗ���
�
�6�9����J���� T��h]��F���9�
�&�_�w�}�����ơ�CF�N��U����u�k�d�]�}�W���Y����`2��rN��U���u�u�u�u�3�3�(���-���U��=N��U���u�<�d����J���K���F�N�� �����u�k�d�t�W���	����^��d��U���u�6�>�h�w�-����s���F�E����u�%�'�!�]�}�W���Y����[�P�����a�
�e�_�w�}�W������F��G1��*��
�d�_�u�w�}�W������F��G1��*��
�%�:�0�]�}�W���Y���F��G1��*��
�0�_�u�w�}�W������T��Q��A݊�g�n�_�u�w��(�������@9��Y��G���8�-�1�%��}�W���	����GF��\��6���
�
�8�9�d�3�(���
����9��O1�����u�2�;�'�4�0����Y���F��sN��U���u�u�u�u���$���<���JǻN��U���<�e����`�W��s���F�S��*����u�k�f�{�}�W���Yӂ��G9��s:��H���g�_�u�u�8�)����Q���F�
��E��u�'�
� �f�n���Y���F��^ �H���'�
� �d�d�-�[���Y�����CN��U���
� �d�f�'�t�}���YӀ��l ��[1����g�&�f�
��<�(���&�����G�����e�g���1�m����&�Ԣ�lU��D1�*ۊ�4�
�&�_�w�}�����ơ�CF�N��U����u�k�d�]�}�W���Y����`2��rN��U���u�u�u�u�3�3�(���-���U��=N��U���u�<�d����J���K���F�N�� �����u�k�d�t�W���	����^��d��U���u�1�;�u�i�;�(���5����G9��h��D���%�y�u�u�w�}����Y����`9��b"��:���d�
� �d�`�-�[���Y�����CN��U���-� ���#�l�(���H�ѓ�O��=N��U���
�<�:�%�d�3�(���K����	F��Z�����8�f�����(���������\�����u�0�0�<�w�<�W�ԜY���F��S�D�ߊu�u�u�u���#���Y���l�N��Uʱ�;�
���w�c�D��Y���F��X��"����h�u�g�]�}�W���Ӌ��NǻN��U���9�u�k�4��1�[���Y�����R��Kʴ�
�&�y�u�w�}�WϺ������h��D���%�y�u�u�w�}����GӁ��l ��X�����u�u�u�u�3�(�W�������F9��1��\�ߠu�u�3�e�$�)����K����9��bZ��U���%�;�;�u�g�o�6����֓�Z��G1����g�g�u�u�0�3�������9F�N��U���h�u�y�u�w�}�Wϐ�4����t#�	N����u�u�u�<�g�
�3���D����l�N��Uʱ� �
���w�c�D���Y����\��Z��]���u�u�u�6�<�`�W�������F�N�����!�h�u�%�%�)�}���Y���W��S����3�
�c�
�g�W�W���Y�Ư�[�P�����c�
�0�_�w�}�W������F��G1��*��
�d�n�_�w�}�(߁�������\��*ۊ�
�`�o�6�:�2��������r%��Q1�����
�g�&�f�9��(�ԜY�ƫ�]��TN�����u�u�u�u��}�I��s���F�y;��&����h�u�y�w�}�W�������d/��N��U��_�u�u�u�w�4�F���=���F��d��U���u�1� �
��	�W���H���F��E�����_�u�u�u�w�4�G��Y����U�� _��E�ߊu�u�u�u�>�l�J�������lW��h����u�u�u�%�8�8�J�������lW��h�����_�u�u�u�w�2���Y����U�� _��G��_�_�_�u�w�p��������]��C��U´�
��3�8�w�;����
������_��[���_�u�u�%������
����l��TN����0�&�4�
�;�t�W�������9F�N��U���}�%�6�>�2�8�Ͽ�Ӈ��P
��
N��D���!�0�_�u�w�}�W���Y���R��D��U��|�!�0�_�w�}�W���Y���F��h-�����i�u�%���)�(���&��ƹF�N��U���9�0�u�u�w�}�W���Y����UF�V�����
�:�<�
�w�}����P�Ƹ�V�N��U���u�u�u�u�w�}����*����Z�V��&���8�_�u�u�w�}�W���Y�Ʃ�WF��NךU���u�u�u�u�9�}��ԜY���F��SN��N���u�0�1�%�8�8��Զs���K��h_��'���:�<�<�;�6���������@��YN�����&�u�x�u�w�-�F߁�����Z��Y1��*���
�'�2�4�$�:�(�������A	��D�����>�_�u�u�2�4�}���Y���Z �V�����#�;�u�;�w�-����D���O��_��U���u�u�u�u�>�}����
���W������u�u�u�u�w�}�WϮ�Hù��E6��^�����
�9�
�'�0�a�W�������l
��^��N���u�u�u�u�w�8��ԜY���F�N��Uʼ�u�}�%�6�9�)���������T��U���;�u�u�u�w�}�W���Y�����F��*���&�
�:�<��}�W���
����@��d:�����3�8�d�|�w�5��ԜY���F�N��U���u�u�u�%�f�����
����]9��h��*���2�i�u�%�4�3��������l�N��U���u�u�u�u�w�8����Q����Z��S
��D���=�;�_�u�w�}�W���Y���F�N����
�0��&�#�2�(�������A��S��*����#�:�<�>�3������ƹF�N��U���u�u�u�u�9�}��ԜY���F�N��Uʰ�1�<�n�_�w�}�W���Y�Ʃ�WF��d��U���u�0�1�<�l�}�Wϻ�Ӗ��P��dװU���x�u�
�e��+��������A��V�����'�6�&�{�z�W�W���&�֓�V��D�����'�2�4�&�0�����CӖ��P�������_�u�u�0�>�W�W���Y�ƥ�N��h��R���;�u�;�u�'�>���Y�����Yd��U���u�u�u�<�w�<�(���Y���O��_��U���u�u�u�u�w�}���&����\��^�����u�h�4�
�8�.�(���K����F�N��U���0�&�_�u�w�}�W���Y���Z �F��*���&�
�:�<��}�W�������]��X��]���6�;�!�9�0�>�F������T9��R��!���d�3�8�e�w�3�Wǿ�&����G9��P��E��4�
�!�'�~�t����Q����\��h�����u�u�
�e��+��������C9��SG��U���;�_�u�u�w�}�W���Y���F��^�����&�!�:�
�%�:�K���&�֓�V��D����u�u�u�u�w�}�W�������U]�N��U���u�u�0�1�>�f�W���Y����]��QUךU���;�u�'�6�$�f�}���Y���C9��h/��%���!�:�
�%�!�9����Y����T��E�����x�_�u�u��l�6�������\��G1�����0�
�&�<�9�-����Y����V��V�����u�u�7�2�9�}�W���Yӏ����T�����!�4�1�4��1�W���^���G��=N��U���u�u�u�3��-����D����F��R ךU���u�u�u�u�w�}�(���8����@��X �����1�%�0�u�j�<�(���
����T��UךU���u�u�u�u�;�8�W���Y���F�N�����4�
�:�&��2����Y�ƭ�l��N���ߊu�u�u�u�w�}�W���Y�ƥ�N��G1�����9�2�6�d�j�<�(���&����l5��D�*���
�e�|�!�2�}�W���Y���F�N��U���u�u�
�d��.��������C9��S1�����h�4�
�:�$�����&��ƹF�N��U���u�u�u�u�;�4�Wǿ�&����Q��^�����u�u�u�u�w�}�W���Y���F���D���&�:�<�<�9�<�(���&����Z�G1�*����&�!�:��-����s���F�N��U���u�u�0�1�>�f�W���Y���F�N�����3�u�u�u�w�}�W�������U]ǻN��U���;�u�3�_�w�}��������@]Ǒ=N��U���%�d�
�7��.����&������^	�����0�&�u�x�w�}���&����\��^�����
�&�<�;�'�2�W�������@N��h��\���u�7�2�;�w�}�W�������C9��\I�����4�1�4�
�;�}�W���^�Ƹ�VǻN��U���u�u�3�}�'�/���^���G��=N��U���u�u�u�u�w��F���
����G��h����u�%�6�;�#�1�D݁�B���F�N��U���0�u�u�u�w�}�W���Yӏ��N��G1�����9�2�6�d�j�<�(���Y����]	��F��*���&�
�:�<��}�W���
����@��d:��ۊ�&�
�|�4�3�u��������\��h^��U���&�4�!�|�w�3�Wǿ�&����G9��P��D��%�d�
�7��.����&����_�N�����u�u�u�u�w�}�W���Y����lW��v�����<�;�%�0�w�`���&����\��^�����u�u�u�u�w�}�W���Y����9F�N��U���u�;�u�3�]�}�W���Y����Z ��N�����%�:�0�&�]�W�W���TӖ��l��R�����
�9�
�'�0�<����Y����V��C�U���%�c�1��%�8�(�������A��V�����'�6�o�%�8�8�ǿ�&����9F����ߊu�u�u�u�1�u����ԃ��]��Y
�����>�h�u�d�~�)��ԜY���F�N��U´�
�&�u�u�f�t����s���F�N��U���%�c�1��%�8�(�������A��S�����;�!�9�2�4�m�}���Y���F�R�����u�u�u�u�w�}�W���Qۇ��P	��C1�����d�h�4�
�2�t����s���F�N��U���u�u�<�u��-��������Z��S�����2�6�0�
��.�Fށ�
����O��_�����u�u�u�u�w�}�W���Y���C9��S:�����
�%�#�1�'�8�W������]��[����_�u�u�u�w�}�W���Y���V
��QN�����2�7�1�`�~�)����Y���F�N��U���u�u�u�u���#���*����C9��S1�����h�%�c�1��/����	����l�N��U���u�u�u�u�w�8�Ϸ�B���F�N��U���u�;�u�3�w�}�W���Y����������u�u�u�;�w�;�}���Y����C��R���ߊu�u�x�%�a�9�'�������V��D��ʥ�:�0�&�u�z�}�WϮ�O����V��T1�����&�<�;�%�8�}�W�������R��[��U���7�2�;�u�w�}�WϷ�Yۇ��P
��R��ʴ�1�4�
�9�w�}�P���Y����9F�N��U���u�3�}�%�%�)�J���^�Ƹ�VǻN��U���u�u�u�u���#���*����A��S�����;�!�9�f��f�W���Y���F��[��U���u�u�u�u�w�}����Qۇ��P	��C1�����d�h�4�
�2�}��������]��[����h�%�c�1��/����	����F��SN�����4�
�:�&��2����Y�ƭ�l��h�����
�!�
�&��t����Q����\��h�����u�u�%�&�6�)�^���Y����l�N��U���u�u�u�u�w�-�A���)����P9��R	��Hʥ�c�1��'�2�f�W���Y���F�N�����3�u�u�u�w�}�W�������U]ǻN��U���;�u�3�_�w�}��������@]Ǒ=N��U���%�m��#�2���������W9��R	�����;�%�:�0�$�}�Z���YӖ��l4��g�� ���
�%�#�1�'�8�(�������A	��N�����&�4�
�9�~�}�Wϼ���ƹF�N�����%�6�>�0�2�)��������XF�I�\ʡ�0�_�u�u�w�}�W����έ�l��S��D���!�0�_�u�w�}�W���Y���C9��e�����9�0�4�
�;�����E�ƭ�l��D�����
�n�u�u�w�}�W�������F�N��U���u�u�<�u��-��������Z��S�����|�u�=�;�w�}�W���Y���F�N�����4�
�:�&��2����Y�ƭ�l��h�����
�!�d�3�:�l�^������F�N��U���u�u�u�u�w�}����+����A6��D�����1�%�0�u�j�<�(���
����T��UךU���u�u�u�u�w�}�W���������D�����c�|�!�0�w�}�W���Y���F�N��U���u�
�
�0��/����&����_��E��I���
�
�0��%�(����	����l�N��U���u�u�u�u�w�8�Ϸ�B���F�N��U���u�;�u�3�w�}�W���Y����������u�u�u�;�w�;�}���Y����C��R���ߊu�u�x�%�o�����)����l��PN�����u�'�6�&�y�p�}���Y����a��R�����%�0�
�&�>�3����Y�Ƽ�\��DF��*���|�u�u�7�0�3�W���Y����UF��G1��Ͱ�0�!�4�1�6�����Y����F��R ךU���u�u�u�u�1�u�������A�C�����u�u�u�u�w�}�W���&����V��[�����u�h�4�
�8�.�(���K����F�N��U���0�&�_�u�w�}�W���Y���Z �F��*���&�
�:�<��}�W�������]��X��]���6�;�!�9�0�>�F������T9��R��!���d�3�8�e�w�3�Wǿ�&����G9��P��E��4�
�!�'�~�t����Q����\��h�����u�u�
�
�2�����
����l��G�����u�u�u�u�w�}�W���Y�����h<��%��� �&�
�'�0�a�W���&����V��[�����u�u�u�u�w�}�W���Y����9F�N��U���u�;�u�3�]�}�W���Y����Z ��N�����%�:�0�&�]�W�W���TӇ��Z��G�����u�x�u�u�'�2����Q����_�N�����;�u�u�u�w�4�Wǿ�&����V��CN��ʴ�
�9�u�u�f�t����s���F�N�����}�4�
�:�$�����&���R��RG�����4�
�:�&��2����Y�ƭ�l��h�����
�!�
�&��t�^Ϫ����F�N��U���u�7�:�
��$����K����lS��R�����
��,� ��o����Iù��l�N��U���u�0�1�<�l�}�W���YӃ����=N��U���u�'�6�&�l�W�W���TӇ��Z��G�����u�x�u�u�'�2����Q����_�N�����;�u�u�u�w�4�Wǿ�&����V��CN��ʴ�
�9�u�u�f�t����s���F�N�����}�4�
�:�$�����&���R��RG�����4�
�:�&��2����Y�ƭ�l��h�����
�!�
�&��t�^Ϫ����F�N��U���u�7�:�
��$����@����lS��R�����
��,� ��d����LĹ��l�N��U���u�0�1�<�l�}�W���YӃ����=N��U���u�'�6�&�l�W�W���TӇ��Z��G�����u�x�u�u�'�2����Q����_�N�����;�u�u�u�w�4�Wǿ�&����V��CN��ʴ�
�9�u�u�f�t����s���F�N�����}�4�
�:�$�����&���R��RG�����4�
�:�&��2����Y�ƭ�l��h�����
�!�
�&��t�^Ϫ����F�N��U���u�3�
����<���	����9��S��&��� ���!�f�����I��ƹF�N��U���u�u�����8���Jƹ��A��]�I��������)�Dځ�&����P��UךU���u�u�u�u�9�}��ԜY���F��SN��N���u�0�1�%�8�8��ԶY���F��D��U���6�&�{�x�]�}�W���������T�����u�0�<�_�w�}�W����έ�l�������;�u�%�6�<�`�P���Y����9F�N��U���u�3�}�}�'�>��������lW������4�1�}�%�4�3��������[��G1�����0�
��&�e�;���P�Ƹ�VǻN��U���u�u�u�u��3��������V��R	��L���h�2�%�3��k�(��s���F�N��U���3�
�:�0�#�/�(��&����_��S����� �d�b�%�l�}�W���Y���F�������;� �
�n�l����L���F��h��9����!�g�
��(�D���	��ƹF�N��U���;�u�3�_�w�}�W����ƥ�l�N��ʥ�:�0�&�_�w�}�Z���
������T��[���_�u�u�'�4�.�Wǿ�&����9F����ߊu�u�u�u�1�u����ԃ��]��Y
�����>�h�r�r�w�5����Y���F���]���%�6�;�!�;�:���DӇ��P�V ��]���6�;�!�9�0�>�F������T9��R��!���f�3�8�g�~�}����Y���F�N��U����-� ���)�Fہ�����F�	��*���d�f�%�n�w�}�W���Y���F��d1�� ����!�d�
�2��F���DӀ��K+��c����
� �d�b�'�f�W���Y���F��Y
���ߊu�u�u�u�9�}��ԜY�Ʃ�WF��X���ߠu�u�x�u�$�4�Ϯ�����F�=N��U���6�&�u�4��1�^���Yӄ��ZǻN��U���3�}�%�6�<�8��������C9��\N��R��u�=�;�u�w�}�W���Yӏ��N��G1�����9�2�6�d�j�<�(���Y������T�����2�6�d�h�6�����
����g9��^�����|�|�!�0�]�}�W���Y���F�Q=��8���,� �
�c�%�:�B��E�ƫ�C9��h_�*��_�u�u�u�w�}�W���Y����F�N�����<�n�u�u�2�9��������9F�C����2�u�'�6�$�s�Z�ԜY�Ƽ�\��DN�����>�_�u�u�2�4�}���Y���Z �V�����#�;�u�;�w�-����D����F��R ךU���u�u�u�u�1�u�_�������l
��^��U���%�6�|�4�3�u��������\��h_��U���&�2�6�0��	��������O�C�����u�u�u�u�w�}�W�������|��]�����a�u�h�2�'�;�(��&����F�N��U���0�1�<�n�w�}�W�������U]ǻN�����'�6�&�n�]�}�W������V��D�����%��
�&�~�2�W���Y����VF��T�����x�u�u�4����������]9��X��U���6�&�u�4������Y����VJ��G1�����1�l�|�u�w�?����Y���F��V������3�8�<�]�}�W���Y���D����&���!�
�&�
�w�c�}���Y���F�N�����}�4�
�:�$�����&���R��RG�����:�}�%�&�0�?���P����[��N��U���u�u�u�u�w�}����*����Z�V��!���g�3�8�d�]�}�W���Y���F�R�����u�u�u�u�w�}�W���Y����`9��ZN�U����
�!�
�$��L���Y���F�N��U���u�3�_�u�w�}�W���Y������d:��؊�&�
�u�k�]�}�W���Y���F�V��&���8�i�u�%���܁�
����9F�N��U���u�=�;�4��	��������[�=N��U���u�u�u�u�w�-�9���
�����d:��ފ�&�
�n�u�w�}�W���Yӑ��]F��h=�����3�8�f�h�w�}�W���Y���F���;���&�u�h�4��	��������l�N��U���u�"�0�u�'��(���&����F�d��U���u�u�u�u�w�<�(������F��h=�����3�8�`�_�w�}�W���Y�ƻ�V��G1��*���
�&�
�u�i�W�W���Y���F�N��*���3�8�i�u�'��(���&����]ǻN��U���u�u�=�;�6��#���N����lP�	NךU���u�u�u�u�w�}����&����[��G1��*���
�&�
�n�w�}�W���Y����[��V��!���m�3�8�b�j�}�W���Y���F�N�����
�&�u�h�6��#���@����l^��N��U���u�u�"�0�w�-�$���ʹ��^9��
P��U���u�u�u�u�w�}����*����Z�V��!���d�
�&�
�l�}�W���Y�����YN��*���&�d�
�&��}�I�ԜY���F�N��Uʴ�
��3�8�k�}����&����l ��h_����u�u�u�u�w�5�Ͽ�&����GW��Q��D���k�_�u�u�w�}�W���Y�ƭ�l(��Q��I���%��
�!��.�(��Y���F�N�����:�=�'�u�i�}�W���Y���F�N�����
�&�u�h�u��/���!����l�N��Uʰ�1�6�&�n�w�}����	����@��=N��U���4�
�:�0�6�.��������@H�d��Uʴ�
�:�0�4�$�:�(�������A	��D�����y�4�
�<��.����&����l ��h_����u�0�<�_�w�}�W������R��X ��*���<�
�u�u�'�>�^Ͽ��έ�l��D�����
�u�u�%�$�:����&����GW��Q��D���|�!�0�u�w�}�W���Y����C9��Y��Hʴ�
�:�&�
�8�4�(��Y���F��[�����u�u�u�u�w�-����Y����C9��Y�����6�e�_�u�w�}�W���Y����9F���U���6�&�n�_�w�}�Z���	����VF��D��U���6�&�{�x�]�}�W�������R��P �����o�%�:�0�$�<�(�������C9��P1������&�d�3�:�m�}���Y����]l�N��Uʼ�u�}�:�}�6�����&����P9��
N��*���'�|�u�;�w�<�(���
����T��N�����<�
�&�$���ށ�
����O��_�����u�u�u�u�w�-����Y����C9��Y�����6�d�_�u�w�}�W������F�N��Uʴ�
�1�0�i�w�-��������Z��d��U���u�0�1�<�l�W�W����Ƽ�\��DUװ���u�x�4�
�2�9�W�������A	��D�X�ߊu�u�%�'�6�$��������\������}�%�6�y�6�����
����g9��_�����e�_�u�u�2�4�}���Y���Z �F��*���&�
�:�<��}�W�������]�V�����
�:�<�
�w�}��������B9��h��D���8�d�|�|�#�8�W���Y���F������,�i�u�%�4�3��������l�N��Uʰ�&�u�u�u�w�}�W�������R��S�����;�!�9�2�4�m�}���Y���V��^����u�;�u�'�4�.�L�ԶY���F��h��*���
�d�u�&�>�3�������KǻN�����2�7�1�d�d�<����&����\��E�����%��
�&�~�}�Wϼ���ƹF�N��U���u�u�%�&�0�?���J�����T�����d�d�h�4������Hӂ��]��G����u�;�u�'�4�.�L�ԶY���F��h��*���
�g�u�&�>�3�������KǻN�����2�7�1�d�`�<����&����\��E�����%��
�&�~�}�Wϼ���ƹF�N��U���u�u�%�&�0�?���N�����T�����d�d�h�4������Kӂ��]��G����u�;�u�'�4�.�L�ԶY���F��h��*���
�f�u�&�>�3�������KǻN�����2�7�1�d�n�<����&����\��E�����%��
�&�~�}�Wϼ���ƹF�N��U���u�u�%�&�0�?���@�����T�����d�d�h�4������Jӂ��]��G����u�;�u�'�4�.�L�ԶY���F��h��*���
�a�u�&�>�3�������KǻN�����2�7�1�d�n�<����&����\��E�����%��
�&�~�}�Wϼ���ƹF�N��U���u�u�%�&�0�?���@�����T�����d�d�h�4������Oӂ��]��G����u�;�u�'�4�.�L�ԶY���F��h��*���
�c�u�&�>�3�������KǻN�����2�7�1�d�f�<����&����\��E�����%��
�&�~�}�Wϼ���ƹF�N��U���u�u�%�&�0�?���H�����T�����d�d�h�4������Nӂ��]�� G����u�;�u�'�4�.�L�ԶY���F��h��*���
�b�u�&�>�3�������KǻN�����2�7�1�d�f�<����&����\��E�����%��
�&�~�}�Wϼ���ƹF�N��U���u�u�%�&�0�?���H�����T�����d�d�h�4������Aӂ��]��G����u�;�u�'�4�.�L�ԶY���F��h��*���
�m�u�&�>�3�������KǻN�����2�7�1�d�g�<����&����\��E�����%��
�&�~�}�Wϼ���ƹF�N��U���u�u�%�&�0�?���I�����T�����d�d�h�4������@ӂ��]��G����u�;�u�'�4�.�L�ԶY���F��h��*���
�m�u�&�>�3�������KǻN�����2�7�1�d�n�<����&����\��E�����%��
�&�~�}�Wϼ���ƹF�N��U���u�u�%�&�0�?���@�����T�����d�d�h�4������H�ƨ�D��_�\�ߊu�u�;�u�%�>���s���K�V�����1�
�e�u�$�4�Ϯ�����F�=N��U���&�2�7�1�e�o��������\������}�%��
�$�t�W�������9F�N��U���u�u�u�%�$�:����K���F��G1�����9�d�d�h�6��$�������\��XN�\�ߊu�u�;�u�%�>���s���K�V�����1�
�b�4�$�:�W�������K��N�����<�
�1�
�`�<����&����\��E�����%��
�&�~�}�Wϼ���ƹF�N��U���u�u�%�&�0�?���Y���R��d1����1�"�!�u�~�`��������_��G�U���0�1�%�:�2�.�}�ԜY�����D�����f�g�4�&�0�}����
���l�N��*���
�1�
�m��.����	����	F��X��´�
��3�8�]�}�W������F�N��U���u�4�
�<��9�(��Y���R��X ��*���
�u�u�%������Y����G	�G�U���0�1�%�:�2�.�}�ԜY�����D�����`�u�&�<�9�-����
���9F������7�1�`�
�$�4��������C��R�����!�'�y�4��4�(�������@��Q��E���
�
��0��>������ƹF��R	�����u�u�u�u�w�}�W���
����W��N�U���%�6�;�!�;�:���DӖ��l��R�����
�9�|�4�3�3��������]��[����h�4�
�<��.����&����U��G�����4�
�:�&��2����Y�ƭ�l��E��\��u�u�0�1�'�2����s���F������7�1�c�u�$�4�Ϯ�����F�=N��U���&�2�7�1�a���������PF��G�����4�
�!�'�{�<�(���&����l5��D�����e�u�
�
�2�����
����l��d��Uʷ�2�;�u�u�w�}�W���Y����C9��P1����u�h�}�:��u��������\��h_��U���&�2�6�0��	��������F��SN�����;�!�9�2�4�m�JϿ�&����GO���U´�
�:�&�
�8�4�(���Y����a��R�����4�
�9�|�l�}�Wϻ�Ӗ��P��dװU���x�u�%�&�0�?���Y����T��E�����x�_�u�u�'�.��������R��P �����o�%�:�0�$�<�(�������C9��P1������&�d�3�:�m�W���I����c	��C��*���#�1�_�u�w�8��ԜY���F�N��Uʴ�
�<�
�1��l�K��������T�����2�6�d�h�6�����
����g9��1����u�;�u�4��2��������F�V�����|�|�4�1��-��������Z��S��*����#�:�<�>�3�������9F���U���6�&�n�_�w�}�Z���	����l��hV����2�u�'�6�$�s�Z�ԜY�ƭ�l��h��*���4�&�2�
�%�>�MϮ�������D�����%�&�2�6�2��#���H����lV�G1�*����&�!�:��-����s���Q��Yd��U���u�u�u�u�w�<�(���&����V�
N�����}�%�6�;�#�1����H����C9��P1������&�d�3�:�m�W���Yۇ��P	��C1�����e�h�4�
�#�/�^������R��X ��*���<�
�u�u��l�6�������\��G1�����_�u�u�;�w�/����B��ƹF�N��*���
�1�
�`�6�.��������@H�d��Uʴ�
�<�
�1��h��������\������}�%�&�4�#�}�(ف�-����V��G1�����
�<�y�%�o�����)����l��A�����<�y�%�d��8�'�������R��[
�����2�u�
�d��.��������C9��S1��*���|�u�u�7�0�3�W���Y���F�N�����2�7�1�l�w�`�_Ǯ�H¹��@6��^�����
�9�
�;�$�:�JϿ�&����G9��P��E���'�}�
�e��+��������C9��S1��*���u�u�%�6�9�)�������\�G1��'���0��9�0�6���������[��G1�����9�2�6�e�w�/�_���&����A5��h�����<�
�<�u�w�-��������Z��N��U´�
�!�'�u�w�-��������Z��G�U���0�1�%�:�2�.�}�ԜY�����D�����
��&�d��.�(���
������T��[���_�u�u�%�$�:����&����GW��Q��L���&�2�
�'�4�g��������C9��P1����e�_�u�u�2�4�}���Y���Z �V�����1�
�m�|�#�8�W���Y���F������6�0�
��$�l�(���&�����T�����2�6�d�_�w�}�W������F�N��U���4�
�<�
�$�,�$����֓�@��R�����:�&�
�:�>��L���Y�������U���u�0�1�%�8�8��Զs���K��G1�����0�
��&�f�����IӇ��Z��G�����u�x�u�u�6�����
����g9��_�����e�4�&�2��/���	����@��G1�����1�d�l�_�w�}����s���F�^�����<�
�1�
�o�t����Y���F�N��U���&�2�6�0��	���&����V�
N��*���&�
�:�<��f�W���Y����_��=N��U���u�u�u�%�$�:����&����GW��Q��D���h�4�
�:�$�����&��ƹF�N�����3�u�u�u�2�9��������9l�N�U���&�2�6�0��	����������^	�����0�&�u�x�w�}��������V��c1��D���8�e�4�&�0�����CӖ��P�������7�1�g�|�w�}�������F���]���&�2�7�1�e�t����Y���F�N��U���&�2�6�0��	��������Z�V�����
�:�<�
�l�}�W���YӃ��VFǻN��U���u�u�%�&�0�>����-����l ��h^��Hʴ�
�:�&�
�8�4�(��Y���F��Y
�����u�u�0�1�'�2����s���F������6�0�
��$�o����HӇ��Z��G�����u�x�u�u�6�����
����g9��1�����4�&�2�
�%�>�MϮ�������D�����d�f�_�u�w�8��ԜY���F��F��*���
�1�
�d�~�)����Y���F�N�����2�6�0�
��.�E������F��h�����:�<�
�n�w�}�W�������9F�N��U���u�%�&�2�4�8�(���
�ԓ�@��R�����:�&�
�:�>��L���Y�������U���u�0�1�%�8�8��Զs���K��G1�����0�
��&�d�;�������]F��X�����x�u�u�4��4�(�������@��Q��G���&�2�
�'�4�g��������C9��P1����b�_�u�u�2�4�}���Y���Z �V�����1�
�g�|�#�8�W���Y���F������6�0�
��$�n����K���R��X ��*���<�
�n�u�w�}�Wϻ�
��ƹF�N��U���%�&�2�6�2��#���J����lT�
N��*���&�
�:�<��f�W���Y����]��QU��U���0�1�%�:�2�.�}�ԜY�����D�����
��&�a�1�0�DϿ�
����C��R��U���u�u�4�
�>�����*����9��Z1�����2�
�'�6�m�-����
ۇ��@��U
��D��_�u�u�0�>�W�W���Y�ƥ�N��h��*���
�f�|�!�2�}�W���Y���F��G1�����0�
��&�c�;���E�ƭ�l��D�����
�n�u�u�w�}����Y���F�N��U���&�2�6�0��	��������Z�V�����
�:�<�
�l�}�W���YӃ����d��Uʰ�1�%�:�0�$�W�}���Y����C9��P1������&�`�3�:�i�����Ƽ�\��D@��X���u�4�
�<��.����&����U��1�����
�'�6�o�'�2��������T9��S1�G�ߊu�u�0�<�]�}�W���Y���R��^	�����e�|�!�0�w�}�W���Y�����D�����
��&�`�1�0�C��Y����\��h�����n�u�u�u�w�8����Y���F�N�����2�6�0�
��.�B������F��h�����:�<�
�n�w�}�W�������U]�N�����%�:�0�&�]�W�W���TӇ��@��T��*���&�c�3�8�b�<����Y����V��C�U���4�
�<�
�$�,�$���Ź��^9��V�����'�6�o�%�8�8�ǿ�&����Q��V����u�0�<�_�w�}�W����έ�l��h��*��|�!�0�u�w�}�W���Y����C9��P1������&�c�3�:�h�K���	����@��X	��*��u�u�u�u�2�.�W���Y���F������6�0�
��$�k����L���R��X ��*���<�
�n�u�w�}�Wϻ�ӏ��l�N��ʥ�:�0�&�_�]�}�W������T9��R��!���b�3�8�c�6�.��������@H�d��Uʴ�
�<�
�&�&��(���&����9��D��*���6�o�%�:�2�.��������W9��GךU���0�<�_�u�w�}�W���Q����Z��S
��A���!�0�u�u�w�}�W���YӇ��@��T��*���&�b�3�8�a�a�W�������l
��^��N���u�u�u�0�$�}�W���Y���F��G1�����0�
��&�`�;���E�ƭ�l��D�����
�n�u�u�w�}�������F�R �����0�&�_�_�w�}�ZϿ�&����P��h=�����3�8�b�4�$�:�W�������K��N�����<�
�&�$���ׁ�
����R��P �����o�%�:�0�$�<�(���&����P��=N��U���<�_�u�u�w�}����	����l��h_�\ʡ�0�u�u�u�w�}�W�������T9��R��!���m�3�8�b�k�}��������\��h_�U���u�u�0�&�w�}�W���Y�����D�����
��&�m�1�0�@��Y����\��h�����n�u�u�u�w�8�Ϸ�B���F��SN�����&�_�_�u�w�p��������V��c1��L���8�m�4�&�0�}����
���l�N��*���
�&�$���)�(���&˹��@��h����%�:�0�&�6���������OǻN�����_�u�u�u�w�;�_���
����W�� _�����u�u�u�u�w�}�WϿ�&����P��h=�����3�8�m�i�w�-��������Z��d��U���u�0�&�u�w�}�W���Y����C9��P1������&�l�3�:�e�K���	����@��X	��*��u�u�u�u�2�9���s���V��G�����_�u�u�7�8��0�������l ��^�����h�}�8�
��(�D���	�ƭ�WF��G1��*��
�g�n�u�w�?����5����G9��h��A���%�u�h�}�:��G���&����CT��Y
����� �d�d�%�~�W�W���*����v%��B��@���3�
�d�
�d�a�W���Y�����h��D���%�u�=�;��2����-����lU��E��@��e�u�u�d�~�8����Y���F��d1�� ����!�d�
�2��F��Y����`9��{+��:���f�
�
�:�>�)����K����Z�Q=��0���� �
�`�e�/���K���F��h��9����!�g�
��(�D���	���l�N��Uʳ�
���g��)�Eց�����l��@��U¦�9�!�%�
�"�n�E���Q���A��N�����u�u�u�u�'�e�%�������@��Y1���ߊu�u��-��	����&�ߓ�F9��1��U��%��&�9�����M����9F�������;� �
�n�4�(���&����U��Z��G��u�!�
�:�>�����ۓ��Z��SF��'���9�
�
� �e�k����Rӓ��Z��SF��*���&�
�#�m�f�t�}���Y����~3�� ����
�;�3��'����A����[�N��U���'�!�g�<�>�>��������F9��1��U���;�}�0�
�:�o����M����V�
N��R���9�0�_�u�w�}�W���&����U��V��F�ߊu�u��-��	�8���HĹ��lW��h�I����;�1�
�2�0�F�������
T��N�������,� ��j����LĹ��Z�Q=��8���g��!�g������I��ƹF��d1�� ����!�d�
�8�4����&����CW�
N��*����,� �
�`�/���M��ƹF�N�����
�a�
�0�6�.��������@H�d��Uʲ�%�3�
�a��8��������\������}�%�6�y�5�2�(��� ���� T��R	��G���4�
�<�
�$�,�$���Ĺ��^9���������!�f��8�(��UӇ��@��T��*���&�m�3�8�`�}��������B9��h��*���
�y�4�
�>�����*����V��D��Yʴ�
�<�
�&�&��(���H����lW�������6�0�
��$�h����M�ƭ�l��h�����
�!�
�&��t�W�������9F�N��U���}�}�%�6�9�)���������T�����}�4�
�:�$�����&���R��^	������
�!�
�$��^ϱ�Yۇ��P	��C1�����d�h�4�
�>�����*����9��Z1�U���}�%�6�;�#�1����H����C9��P1������&�l�3�:�e�W���Qۇ��P	��C1�����d�h�4�
�>�����*����9��Z1�U���u�:�}�7�8��0�������l��h[�U���%�6�;�!�;�l�G���Y���]	���������!�f��8�(��Y�ƭ�l��D��ۊ�|�u�;�u�6�����&����P9��
N��*���
�&�$���)�(���&���\������!�9�2�6�f�`��������V��c1��Dڊ�&�
�|�4�3�3��������2��B��L���2�`�e�h�6�����&����O���]´�
�:�&�
�8�4�(���Y����Z��D��&���!�d�3�8�f�t�������Q	��h�����
�l�'�2�b�m�JϿ�&����G9��1�\���|�!�0�u�w�}�W���Y����A��B1�B���u�h�4�
�8�.�(�������9F�N��U���0�_�u�u�w�}�W�������lW��h��I���%�6�;�!�;�:���s���F�R ����_�u�u�;�w�/����B��ƹF�N�����
�a�
�%�8�8�����Ƽ�\��D@��X���u�2�%�3��i�(�������@��Y1�����u�'�6�&��2����-����lU��E��@��u�%�&�2�4�8�(���
�ѓ�@��N������,� �
�n�/���I�ƭ�l��h�����
�!�
�&��q��������V��c1��@���8�a�_�u�w�8��ԜY���F��F�����;�!�9�2�4�l�JϿ�&����P��h=�����3�8�c�|�#�8�W���Y���F�	��*���d�b�:�6�3�}�JϿ�&����G9��1����u�u�u�9�>�}�_���	����@��X	��*���u�%�&�2�4�8�(���
�ӓ�@��N��ʻ�!�}�:�9�/�	�8���J����T9��N�����:�&�
�#��t�^ϱ�Y�έ�l��D�����
�u�u�%�$�:����&����G_��D��\ʴ�1�;�!�}�8�1����6����
9��P1�E��4�
�:�&��+�(���P����[��=N��U���u�u�u�'��(�F�������VF������!�9�g�e�]�}�W���Y����l�N��U���u�2�%�3��i�(������F��oL�U���u�u�0�1�>�f�}���Y����C��R���ߊu�u�x�2�'�;�(��&����@��YN�����&�u�x�u�w�:����&����CV��D�����:�u�u�'�4�.�_�������J)��h_�����`�b�u��/��#�������A��_�U���&�2�6�0��	��������F��h=��0��� �
�`�g�%�:�B��Y����Z��D��&���!�
�&�
�{�<�(���&����l5��D�����a�_�u�u�2�4�}���Y���Z ������!�9�2�6�f�`��������V��c1��L���8�m�|�!�2�}�W���Y���F��E�� ��b�%�u�h�1��2���-���� S��h��*��n�u�u�u�w�8����Qۇ��P	��C1�����d�h�4�
�>�����*����9��Z1�\ʡ�0�u�u�u�w�}�W�������F9�� 1��U��3�
���.�(�(�������Q��N��U���0�&�3�}�6�����&����P9��
N��*���
�&�$���)�(���&���G��d��U���u�u�u�2�'�;�(��&���F��h��9��� �
�b�'�0�h�C�ԜY���F��D��U���u�u�u�u�0�-����MĹ��Z�6��-���������/���!����k>��UךU���u�u�;�u�1�}�W�������A	��D����u�x�u�'��(�F���	�ƭ�@�������{�x�_�u�w�/�(���H�ѓ�9��D��*���6�o�%�:�2�.����<����p-��C��*���e�u�%�&�0�>����-����l ��hX����<�
�&�$���ց�
������D�����
��&�`�1�0�C�ԜY�Ʈ�T��N��U���<�u�}�%�4�3��������[��G1�����0�
��&�n�;���PӒ��]FǻN��U���u�u�'�
�"�l�@���Y����C9��Y����
�e�e�e�g�W�W���Y�Ʃ�@��F��*���&�
�:�<��}�W���
����@��d:��݊�&�
�|�u�?�3�}���Y���F�P�����a�
�d�i�w��1���;����F��C1�*��u�u�u�u�2�.��������]��[����h�4�
�<��.����&����U��G�����u�u�u�u�w�}�WϹ�	����R��G_��Hʴ�
�:�&�
�!�o�4��I����9F�N��U���0�_�u�u�w�}�W�������lW��h�I���������/���!����k>��o6��-���n�u�u�u�w�8�Ϸ�B���F��SN�����&�_�_�u�w�p�������� 9�������%�:�0�&�w�p�W�������F9��1��*���<�;�%�:�w�}����
�Ϊ�l��R1�����d�
�0�
�n�q��������V��c1��F���8�g�u��/�����&�Փ�V��[������,� ��k����L���R��^	������
�!�e�1�0�N���	����l��F1��*���d�3�8�d�~�}�Wϼ���ƹF�N�����4�
�:�&��2����Y�ƭ�l��h�����
�!�d�3�:�l�^������F�N��U���2�%�3�
�b��G��Y����~3��N!��*���'�2�`�e�]�}�W���Y����UF�V�����
�:�<�
�w�}��������B9��h��E���8�l�|�!�2�}�W���Y���F��E�� ��f�%�u�h�1��$���6���� 9��P1�@�ߊu�u�u�u�;�4�W���	����@��X	��*���u�%�&�2�4�8�(���
�Փ�@��G�����_�u�u�u�w�}�W���&����U��N�U���;�1�
�0�:�l�C�������l�N��Uʰ�&�u�u�u�w�}�W�������F9��1��U��w������/���!����k>��o6��-���w�_�u�u�w�}������ƹF��Y
�����&�n�_�u�w�p�W���&����U��N�����u�'�6�&�y�p�}���Y����U��]��D���&�2�
�'�4�g��������lP��c>��&���<�
�<�y�'�e�%�������@��Y1�����%�&�2�6�2��#���J����lT�V�����&�$��
�#�m����@�ƭ�l��h�����
�!�d�3�:�l�^���Yӄ��ZǻN��U���3�}�4�
�8�.�(�������F��h��*���$��
�!�f�;���P�Ƹ�V�N��U���u�u�2�%�1��B܁�H���R��X ��*���g�a��e��f�W���Y����_��F�����;�!�9�2�4�l�JϿ�&����P��h=����
�&�
�|�w�5��ԜY���F�N�����
�`�
�d�k�}�(ف�-����V��Y1���ߊu�u�u�u�;�4�W���	����@��X	��*���u�%�&�2�4�8�(���
�Փ�@��G�����_�u�u�u�w�}�W���&����U��N�U���
�0��'�"�.�(���
����F�N�����u�u�u�u�w�}�WϹ�	����S��G_��H���������/���!����k>��o6��-���_�u�u�u�w�3�W���Y����������n�_�u�u�z�}��������l��V�����'�6�&�{�z�W�W�������lW��h�����2�
�'�6�m�-����
ۇ��@��T��*���&�d�3�8�g�}����UӇ��@��U
��L���4�
�<�
�$�,�$�������^9��=N��U���<�_�u�u�w�}����Q����\��h�����u�u�%�6�~�<����Q����\��h�����u�u�%�&�0�>����-����l ��h^�����;�!�4�
�>�����L����AF��G1�����9�2�6�d�j�<�(���&����l5��D�����d�|�|�!�2�}�W���Y���F��E�� ��f�6�u�h�6�����&����P9��=N��U���u�9�0�_�w�}�W���Y�ƫ�C9��h_�*���i�u�%�6�9�)��������F�N�����<�n�_�u�w�3�W�������9l�N�����
�c�
�e�k�}�(���+����@��X �����2�_�u�u�z�}��������l��V�����'�6�&�{�z�W�W�������lW��h�����2�
�'�6�m�-����
ۇ��@��T��*���&�d�3�8�g�}����UӇ��@��U
��L���4�
�<�
�$�,�$�������^9��=N��U���<�_�u�u�w�}����Q����\��h�����u�u�%�6�~�<����Q����\��h�����u�u�%�&�0�>����-����l ��h^�����;�!�4�
�>�����L����AF��G1�����9�2�6�d�j�<�(���&����l5��D�����d�|�|�!�2�}�W���Y���F��E�� ��b�6�u�h�6�����&����P9��=N��U���u�9�0�_�w�}�W���Y�ƫ�C9��h_�*���i�u�%�6�9�)��������F�N�����<�n�_�u�w�3�W�������9l�N�����
�c�
�e�k�}�(���8����@��X �����2�_�u�u�z�}��������l	��X
�����2�u�'�6�$�s�Z�ԜY�ƫ�C9��h_�*���:�0�4�&�0�����CӖ��P�������6�0�
��$�i����J�ƭ�l��h�����
�!�
�&��t�W�������9F�N��U���}�4�
�:�$�����&���R��^	������
�!�
�$��^������F�N��U���2�%�3�
�`��������R��X ��*���
�n�u�u�w�}��������C9��Y�����6�d�h�4��4�(�������@��Q��F���!�0�u�u�w�}�W���YӁ��l ��Y�����1�u�h�4��2����ƹ��9F�N��U���0�_�u�u�w�}�W�������lW��h�����i�u����f�W���Y����]��QU��U���0�1�%�:�2�.�}�ԜY�����h��D���%�u�&�<�9�-����
���9F�	��*���d�d�%�
�$�4��������C��R�������,� ��j����L���R��^	������
�!�
�$��[ϸ�&����p2��C1�*؊�0�
�f�y�6�����
����g9��1����_�u�u�0�>�W�W���Y�ƥ�N��G1�����9�2�6�d�j�<�(���&����l5��D�����b�|�!�0�w�}�W���Y�����h��D���%�u�h�3���2�������lT��R	��F��u�u�u�u�2�.��������]��[����h�4�
�<��.����&����U��G�����u�u�u�u�w�}�WϹ�	����Q��G^��Hʳ�
���,�"��@�������l�N��Uʰ�&�u�u�u�w�}�W�������F9��1��U��w������/���!����k>��o6��-���w�_�u�u�w�}������ƹF��Y
�����&�n�_�u�w�p�W���&����W��N�����u�'�6�&�y�p�}���Y����U�� _��D���&�2�
�'�4�g��������C9��P1������&�a�3�:�n�W���
����@��d:��Ҋ�&�
�|�u�w�?����Y���F��QN�����:�&�
�:�>��W���	����l��F1��*���
�&�
�|�w�5��ԜY���F�N�����
�b�
�d�k�}��������EU��u(�E��n�u�u�u�w�8����Qۇ��P	��C1�����d�h�4�
�>�����*����9��Z1�\ʡ�0�u�u�u�w�}�W�������F9��1��U��4�
�:�&��+�E���A����]ǻN��U���9�0�_�u�w�}�W���Y����U�� _��D��u������/���!����k>��o6��-����n�u�u�w�}�������F�R �����0�&�_�u�w�1����H����_��G_��Hʥ��9�
�
�"�l�@���Q���W��X����n�u�u�9�4�����Aù��Z�G1��؊�
� �d�b�'�u�GϺ�����U�=N��U���9�&�
� �c�d����D������YN�����
� �a�`�'�}�W�������l
��h(��U���0�w�w�_�w�}����
���� ^��G\��H���w�"�0�u�#�-�N���&����CR������!�9�m��~�8����H��ƹF��X��ۊ� �a�`�%�w�`�U���������h_�����f�
�d�h�6�����&����lV�R��U��n�u�u�;�#�5�(���J�ޓ�F�L�U���;�}�8�
�b�;�(��&�����T�����g�
�|�0�$�}�G��Y����lV��1�����m�
�f�i�w�}�W���YӇ��P	��C1��Gي�u�=�;�}�:����K����O�I�\ʰ�&�u�u�u�w�}����/�ד�F9��1��N���u�%�e��3�8�$���E�ƫ�C9��h_�*��_�u�u�x�w��(���)����P9��h��U���<�;�%�:�2�.�W��Y����lV��V
�����
�%�#�1�6�.���������T��]���6�y�4�
�>�����*����W��D��E�ߊu�u�0�<�]�}�W���Y���N��h�����:�<�
�u�w�-�������R��X ��*���<�
�u�u�'�.��������l��1����|�|�!�0�w�}�W���Y�����h<��%���0�
�%�#�3�a�W�������l
��^��N���u�u�u�0�$�}�W���Y���F��h^�����'�0�
�%�!�9�K���	����@��X	��*��u�u�u�u�2�9���s���V��G�����_�_�u�u�z�-�F߁�����Z��Y1��*���
�;�&�2�6�.��������@H�d��Uʥ�d�
�0��$�)����	����l��D�����2�
�'�6�m�-����
ۖ��9��A>�����;�4�
�9�{�-�F߁�����Z��Y1��*���
�'�2�_�w�}����s���F�^��]���6�;�!�9�0�>�F��	����a��X�����4�
�9�|�w�5��ԜY���F�N��Dڊ�0��&�!�8���������@��S��*����#�:�<�>�3������ƹF�N�����_�u�u�u�w�}�W���I����c	��C��*���#�1�<�
�>�}�JϮ�Hù��E6��^�����
�9�
�'�0�W�W���Y�Ʃ�WF��NךU���;�u�'�6�$�f�}���Y���C9��h<��%���!�:�
�;�$�:�����Ƽ�\��D@��X���u�%�d�
�2���������l��h�����%�:�u�u�%�>����&�֓�V��D�����%�d�
�0��.����&����F��^�����&�!�:�
�'�+��ԜY�Ʈ�T��N��U���<�u�}�%�4�3��������[��h_��'���:�<�<�;�6�����Y����l�N��U���u�%�d�
�2���������l��R����
�0��&�#�2�L���Y�����RNךU���u�u�u�u��m�%�������\��Y1����u�
�e��!�2��������T]ǻN��U���;�u�3�u�w�}����	����@��=d��U���u�
�d��$�2��������E
��^ �����&�<�;�%�8�8����T�����1�����<�<�;�4��1�(���
����@��Y1�����u�'�6�&���F���
����G��h�����u�
�d��$�2��������E
��G��\���u�7�2�;�w�}�W������R��X ��*���<�
�u�u��l�6�������\��G1�����!�0�u�u�w�}�W���YӖ��9��D>�����;�4�
�9��3����E�Ƽ�W��U�����:�
�%�#�3�W�W���Y�Ʃ�@�N��U���u�u�%�d��?�'�������R��[
�����2�i�u�
�f���������l��A�����n�u�u�u�w�8�Ϸ�B���F��SN�����&�_�_�u�w�p���&����\��^�����<�u�&�<�9�-����
���9F���D���&�:�<�<�9�4�(���&����T��E��Oʥ�:�0�&�%�f�����
����]J��h_��4���:�<�<�;�'�8�[Ϯ�H¹��@6��^�����
�9�|�u�w�?����Y���F��QN�����:�&�
�:�>��W���&�ד�Q��D�����%�#�1�|�#�8�W���Y���F���D���&�:�<�<�9�4�(���Y����lW��v�����<�;�_�u�w�}�W������F�N��Uʥ�d�
�7��$�)��������Z�G1�*����&�!�:��/��ԜY���F��SN��N�ߊu�u�;�u�%�>���s���C9��c����u�u�u�u�w�:����&����CT��_��]���9�-���#�n�(���&����O�I�\ʰ�&�u�u�u�w�}����<����|��[��*���
�f�n�_�w�}�ZϮ�H����G��G1��ʴ�&�2�u�'�4�.�Y��s���C9��c�����
�9�
�&�>�3����Y�Ƽ�\��DF��*���u�%�&�2�4�8�(���
����U��^��U���7�2�;�u�w�}�WϷ�Y����C9��Y�����6�d�h�4��8�W���Yۇ��P	��C1�����d�h�4�
�>�����*����W��D��E���u�=�;�_�w�}�W���Y�Ƽ�9��R�����9�u�h�4��2��������]ǻN��U���9�0�_�u�w�}�W���Y����g��V1��*���u�h�4�
�8�.�(�������9F�N��U���u�3�u�u�w�8�Ϯ�����lǻN��*؊�0��'�0�w�`����4����|��X�����`�n�_�u�w�p����+����A5��h�����4�&�2�u�%�>���T���F��1������6�4�
�;���������PF��G�����4�
�0�u�'�.��������l��1����|�u�u�7�0�3�W���Y����UF������!�9�2�6�f�`�����ƭ�WF��G1�����9�2�6�d�j�<�(���&����l5��D�*���
�e�|�u�?�3�}���Y���F�G1��'���0��6�4��1�W������]��[����_�u�u�u�w�1��ԜY���F�N��G���#�0��6�6�����DӇ��P	��C1�����e�_�u�u�w�}������ƹF��Y
�����&�n�_�u�w��(�������\��S��&��� ���!�f�����I��ƓF�C��*ي�0�:� �<�9�����Ӈ��Z��G�����u�x�u�u�'�n�%�������]��G1�����&�2�
�'�4�g��������C9��N��*���
�&�$���)�F�������9F����ߊu�u�u�u�1�u�_�������l
��^��U���%�6�|�4�3�u��������\��h_��U���&�2�6�0��	���&����V�N�����u�u�u�u�w�}����+����F��Y�����1�i�u�%�4�3��������l�N��Uʰ�&�u�u�u�w�}�W���	�Փ�V��B�����%�#�1�i�w�-��������Z��d��U���u�0�1�<�l�W�W����Ƽ�\��DUװ���u�x�%�c�3�����&����_��Y1��ʴ�&�2�u�'�4�.�Y��s���C9��S:�����
�%�#�1�>�����
����l��TN����0�&�%�c�3�����&����_�G1�����'�0�
�%�!�9����P�����^ ךU���u�u�3�}�6�����&����P9��
N��C����'�0�
�'�+��������9F�N��U���u�
�
��2�����&����Z��^	��Hʥ�c�1��'�2��������F�N�����u�u�u�u�w�}��������`��V�����;�&�2�i�w��(�������l��A�����n�u�u�u�w�8�Ϸ�B���F��SN�����&�_�_�u�w�p��������`��^ �����&�<�;�%�8�8����T�����h
�����6�<�
�<��.����	����	F��X��¥�c�1��'�2�q��������`��G��Yʥ�c�1��'�2��������F��P��U���u�u�<�u��-��������Z��S��*܊��0��6�6�����Y����l�N��U���u�%�c�1��/��������Z�G1�����'�0�n�u�w�}�Wϻ�
��ƹF�N��U���
�
��0��>���������h
�����6�%�0�n�w�}�W�������U]�N�����%�:�0�&�]�W�W���TӖ��l4��g�� ���
�%�#�1�>�����
������T��[���_�u�u�
��8�'�������R��[
�����2�4�&�2��/���	����@��hV�����'� �&�
�'�+����&˹��E6��g�����
�9�
�'�0�W�W�������F�N�����}�%�6�;�#�1����H����l^��R�����&�
�%�#�3�t����Y���F�N��U���
�0��'�"�.�(�������]9��PN�U���
�0��'�"�.�(�������F�N�����u�u�u�u�w�}�WϮ�A����c��B��*���#�1�<�
�>�}�JϮ�A����c��B��*���#�1�%�0�l�}�W���YӃ����d��Uʰ�1�%�:�0�$�W�}���Y����l^��R�����&�
�;�&�0�<����Y����V��C�U���%�m��#�2���������T9��D��*���6�o�%�:�2�.����+����A6��D�����#�0��;�8����UӖ��l4��g�� ���
�%�#�1�]�}�W������F�N��U���%�6�;�!�;�:���DӖ��l4��g�� ���
�%�#�1�~�)����Y���F�N��*Ҋ�0��'� �$��������C9��e�����9�0�_�u�w�}�W������F�N��Uʥ�m��#�0��1����&����[��hV�����'� �&�
�%�:�}���Y���V��^����u�;�u�'�4�.�L�ԜY�Ƽ�a��[��*���f�a�%�u�j�u�(���K����F9�� 1��]��1�"�!�u�f�}�W���&¹��lU��h�N���u�%��&�;��(���K�Г� F�F��*���&�
�#�e�g�{����/����^��GZ����u�
�4�g�$�;�(��&���F��1������9�0�<��4�L���YӔ��lT��h�����6�&�
� �e�m����D���F�N��*���&�
�#�`�b�m� ���Yے��l^��h�� ��e�%�}�|�j�z�P������F�N�����:�&�
�#�b�l�G�ԜY�ƾ�G9��^1��*��
�f�i�u�w�}�W�������]��[�*��e�"�0�u�#�-�O�������V��G\��\��r�r�u�9�2�W�W���Y�ƭ�l��D�����a�e�n�u�w�.����	¹��lT��h�I���!�%�<�<�1��Nہ�KӞ����T�����d�d�n�u�w�.����	����lT��h�I���!�%�<�<�`�;�(��&����]��R�����3�
�f�
�e�f�W���
����^��Q��Aڊ�g�i�u�d�w�5����*����2��x��Gӊ�;�3��%��(�E���	���R��X ��*���`�a�e�|�2�.�W��B�����h��B���
�a�
�g�k�}�F������U5��z;��G���!�g�
�;�1�	��������l��
N��*���&�
�#�`�c�m�W�������l�N�����%�
� �f�e�-�W��Q����G��h��F���%�u�'�&�;�)�؁�����l��d��Uʦ�9�!�%�3��o�(��E��ƹF�N�����
�
� �g�a�-�W����θ�C9��^1��*��
�g�e�u�w�l�^ϻ�
��ƹF�N�����;�!�9�d��m�L���YӒ��lW��Q��@ۊ�g�i�u�;�#�5�F���&����CT��EN�����d�3�
�f��o�L���YӒ��lW��Q��Eފ�d�i�u��/��#ݰ�����l��R��#���3�
�c�
�e�e�Z������\F��d��Uʡ�%�d�
� �d�e����DӀ��K+��c����
�:�<�!�1��Aځ�H����F��S�����|�_�u�u�:��A���&����CW�
N��*����� �
�b�o��������lR��h�G���u�u�:�;�8�m�L���YӒ��lW��B1�C���u�h�}�8�����A����F��_�*ۊ� �g�m�%�~�W�W�������U��X��F��u�u�u�u�w�<�(���
����9�������8�
�
� �e�m����P���A�R��U���u�u�u�4��2����˹��9F���*ފ� �f�a�%�w�`�_�������F9��1��U���;�!�=�
�"�n�E���P���F��G1�����b�
�g�i�w�l�W����ο�T��������;� �
�n�4�(���&����U��Z��G���u�<�;�1�6�����&����l ��N�����e�n�u�u�#�-�A���&����CT�
N��Wʢ�0�u�&�2�2�u�$���,����|��W�����%��d�3��k�(��Y�ƿ�T�������!�9�d�
�~�}����[����F�C��B���
�g�
�a�k�}�$���5����F��1�����;�
� �a�e�-�_������\F��UךU���8�
�
� �d�e����D���F�N�����3�
�l�
�d�*��������F9��1��]���h�r�r�u�;�8�}���Y���G��\�� ��a�%�n�u�w�)��������F9��1��U��w�w�"�0�w�1����H����_��G_��U���6�;�!�9�e��^ϻ�
���]ǻN�����
� �f�m�'�}�Jϸ�&����g��C1�*���<�!�3�
�a��F��Y����G	�G�U���!�%�3�
�o��E��Yے��lS��B1�E���u�'�!�%�a�;�(��&���9F���*���
�
� �g�c�-�W��[����[����*��� �d�e�%�w�}��������E^��qG�����w�w�_�u�w�0�(���&����
R��N�U��u�=�;�}�8��(���H�֓�F�V�����
�#�
�|�2�.�W��B������V�