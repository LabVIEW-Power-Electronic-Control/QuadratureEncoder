-- � 2012 National Instruments Corporation.
encrypted

�U��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D���[�
d�U���0�2�;�'�#�9��������2��&��U���<�=��#�;�����
����A	��tB��^���;�u�,�!�:�W�Zψ�����	F��Z�����%�'�2�#�u�^��H�Ɣ�_��'��[ʔ�9�'�2�!�w�8�������l�S��H��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D���l��^�����0�0�_�&�w�8��������Z��X����_�0�!�!�w�m�E���=����l ��[1����g�&�f�
��<�(���Y��ƹF��R �����_�u�u�u�w��W���Y�����R	��U��d�_�u�u�w�}�"���-����\��Y�����h�d�_�u�w�}�W���I����g.������u�h�f�n�w�}�W�������d/��N����2�'�o�u�e�W�W���Y�ƨ�F��~*��U���;�0�0�u�j�n�}���Y��ƹF��X��]���u�u�u�1�9�}�W���Y����_	��T1�����}�<�e����FϺ�����O��N��U���1�;�u�u�9�}��������E��X��������d�3�*����P���F�N�� ���u� �u�!��2����������C1��1���d�1�"�!�w�t�W���P���WF��C��N���'�=�!�6�"�8����Y����U��v-�����3� �
�g�$�n����K�ד�R��D�����u�x�x�x�z�p�Z��T���K��X�����u�x�x�x�z�p�Z��T���l�N�����0�!�8�f���6���&����^��1�����%�f�u�&�w�}�W���	����l�N��U���u�&�4�<���������F��^ �����9�2�6�_�w�}�W���Y�ƿ�R��h�����u�u�u�u�w�3�W���&����P9��T��]��1�"�!�u�~�W�W���Y���F��V��*���#�9�1�u�w�}�W���Y����_	��TUךU���u�u�u�u��%��������F�N��U���u�!�
�:�>���������W	��C��\�ߊu�u�u�u�w�}�(���
����F
��C�����u� �u�!��2���Y���F�N��*���&�'�&�9��9����CӉ����h�����0�!�'�f�w�2����I���F�N����u�;�u�:�'�3���Y���K�C�X���x�x�x�x�w�2��������K�C�X���x�x�x�x�w�}�����ƭ�G��^
��U���
�:�<�n�w�}�����ƭ�G��VN��U���
�:�<�
�2�)���Y����G	�UךU���<�;�9�7�#�<����Y����_	��TUךU���<�;�9�7�#�<����Y����_	��T1�����}�d�1�"�#�}�^�ԜY�ƿ�T�������1�o�&�1�;�:��ԜY�ƿ�T�������u�o�&�1�;�:�������� W��X����n�7�2�;�w�}�Z��T���K�C�X���u�;�!�;�>�)����T���K�C�X���u�u�8�f���6���&����^��1�����%�f�
�u�w�2�����ơ� T��t*��*ڊ�%�3� �
��<�(���&��ƹF��X�����}�u�u�u�w�.����&����R
��N��U��u�
�#�9�3�W�W���Y�ƿ�R��h�����u�u�u�u�i�<�������F�N�����
�
�#�9�3�}�W���Gӄ��E��SBךU���u�u�
�-�$�?�������F�	N�����4�_�u�u�w�}�(���
����F
��C�����k�'�!�4�>�q�W���Y����l��D1�����
�1�!�u�j�}�(������F�=d��U���x�x�x�x�z�p�Z��T����@��Y�����x�x�x�x�z�p�Z��T���F��C�����h�r�r�_�w�}�(������F��^ ��"����d�1�"�#�}�W���^���D��F����h�}�1�;���#��Y����G	�S�R��|�u�'�}�>�m�J�������d/��C����!�u�u�k�p�z�^�������Z��=N��U���#�9�1�i�w�l�L���Yӄ��W��N�U±�;�
���z�}�������F�G�����}�1�;�u�w�}����.����W��X����h�u��|�w�2�WǺ����F��Y_��<���x�u�:�;�8�m�J���,�����RN����u�u�1� �w�}�W������G��=��U���=�!�6� �2�W