-- � 2012 National Instruments Corporation.
encrypted

�U��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D���[�
d�U���0�2�;�'�#�9��������2��&��U���<�=��#�;�����
����A	��tB��^���;�u�,�!�:�W�Zψ�����	F��Z�����%�'�2�#�u�^��H�Ɣ�_��'��[ʔ�9�'�2�!�w�8�������l�S��H��h�h�h�h�j�`�J��D���[�
S��H��h�h�h�h�j�`�J��D���l��^�����0�0�_�&�w�8��������Z��X����_�0�!�!�w�m�E���=����l��X��Fػ�
�g�g�<�]�}�W�������l�N��Uʜ�u�u�u�u�w�}��������U��N��U��������}�W�������	[�d��U���u�1�;�
��	�W�������AF��]����u�u�u�:�#�
�3���Cӏ��V��T��F�ߊu�u�n�u�w�-����s���F�T��U��<�u�&�1�;�:��ԜY���F��D��Oʼ�u�&�1�9�0�>�}���Y���P�N����&�1�9�2�4�W�W���Y�ƨ�]V�N��Uʦ�1�9�2�6�!�>�����֓�z"��_�����:�e�n�u�w�}�WϺ����	����*���<�
�0�!�%�9����0����F��@ ��U���u�u�|�_�9�}���� ����A��C�� ���4�6�u�3�:�n�5���8����@��Q��G���f�
�u�&�w�}�Z��T���K�C�X���u�:�%�;�9�}�Z��T���K�C�X���u�u�6�8�8�8�ϳ�J����w'��1��*���:�%�e�;��.�(�����F�N�����_�u�u�u�w�}�W�������l��[��U���u�u�;�u�#�����B���F�N��U���-�&�4�!�6�<�W���Y����]F��C
�����
�0�!�'�d�}�������9F�N��U���u�
�-�&�%�.��������\��B�����:�<�n�u�w�}�W���YӋ��K��E�����1�!�u�o�8�)��������l��C��F���:�;�:�e�]�}�W���Y��ƹF��Y
�����;�;�n�u�w�p�Z��T���K�C�X���:�4�u�<�9�1�Z��T���K�C�X���u�&�2�4�w���������@��[���ߊu�u�<�;�;�<���������h�����0�!�'�f�w�2����I��ƹF��^	��ʧ�!�4�<�u�m�.��������F�D�����
�1�!�u�w�}��������E��X��Dʱ�"�!�u�|�]�}�W�������Z��U��U���!�
�:�<��8��������d/��C����!�u�|�_�2�4�}���Y���K�C�X���x�x�x��$�<�������K�C�X���x�x�_�u�w�m�E���=����l��D�����
�:�1�%�d��W�������V��Z^�7����
�
�%�$�)����&����@��d��Uʥ�'�u�4�u�]�}�W���Y����Z��h�����u�u�u�k�6�)����U���F������4�!�4�4�w�}�W��Y����R��=N��U���u�
�-�&�%�.��������[�E1�����y�u�u�u�w�0����&����_��S��U��u�
�1�!�]�}�W��s���K�C�X���x�x�x�x�z���������K�C�X���x�x�x�x�]�}�W�������Z�_�����u�
�1�!�w�a�WǺ�ù��w2��N�����u�u�k�r�p�}����Qۂ��9��Q_��U���<�e����l��������X�oI��Uʺ�u�1�;�
�"�l�J�������d/��C����!�u�u�k�p�z�^�������Z��U��N���u�1� �u�w�}�JϬ�����lǻN��X���x�x�x�x�z�p�Z��Y����GF��Q��U���x�x�x�x�z�p�Z��Y����A	��D�����u�0�<�_�w�}�W���Ӆ����Y�����9�u�u�d�w�5����Y���F������u�d�u�=�9�}�W���Y���F�
��E���3�u�h�1�9�f�W���Y���F��Y
���ߊu�u�u�u�9�}��ԜY�Ʃ�WF��X���ߠ0�1�4�6�>�8����B�